`timescale 1ns / 1ps
/*******************************************************************************
Company        : AEgis Technologies
Engineer       : John Zartman

Create Date    :
Design Name    :
Module Name    : MODULE_NAME
Project Name   :
Target Devices : Zedboard
Tool Versions  : Vivado 2019.1

Description:

Dependencies:

Additional Comments:

*******************************************************************************/

module MODULE_NAME #(
  parameter
) (
  input wire
  output reg
);

endmodule

